library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

ENTITY binaryToBCD is

	port( input: in std_logic_vector(7 downto 0);
			d1, d2: out std_logic_vector(3 downto 0)
	);
	
end ENTITY;

architecture behv of binaryToBCD is


	begin

		process(input)
		
			begin
			
								CASE input IS
    when "00000000" => d1 <= "0000"; d2 <= "0000"; -- 0
    when "00000001" => d1 <= "0001"; d2 <= "0000"; -- 1
    when "00000010" => d1 <= "0010"; d2 <= "0000"; -- 2
    when "00000011" => d1 <= "0011"; d2 <= "0000"; -- 3
    when "00000100" => d1 <= "0100"; d2 <= "0000"; -- 4
    when "00000101" => d1 <= "0101"; d2 <= "0000"; -- 5
    when "00000110" => d1 <= "0110"; d2 <= "0000"; -- 6
    when "00000111" => d1 <= "0111"; d2 <= "0000"; -- 7
    when "00001000" => d1 <= "1000"; d2 <= "0000"; -- 8
    when "00001001" => d1 <= "1001"; d2 <= "0000"; -- 9
    when "00001010" => d1 <= "0000"; d2 <= "0001"; -- 10
    when "00001011" => d1 <= "0001"; d2 <= "0001"; -- 11
    when "00001100" => d1 <= "0010"; d2 <= "0001"; -- 12
    when "00001101" => d1 <= "0011"; d2 <= "0001"; -- 13
    when "00001110" => d1 <= "0100"; d2 <= "0001"; -- 14
    when "00001111" => d1 <= "0101"; d2 <= "0001"; -- 15
    when "00010000" => d1 <= "0110"; d2 <= "0001"; -- 16
    when "00010001" => d1 <= "0111"; d2 <= "0001"; -- 17
    when "00010010" => d1 <= "1000"; d2 <= "0001"; -- 18
    when "00010011" => d1 <= "1001"; d2 <= "0001"; -- 19
    when "00010100" => d1 <= "0000"; d2 <= "0010"; -- 20
    when "00010101" => d1 <= "0001"; d2 <= "0010"; -- 21
    when "00010110" => d1 <= "0010"; d2 <= "0010"; -- 22
    when "00010111" => d1 <= "0011"; d2 <= "0010"; -- 23
    when "00011000" => d1 <= "0100"; d2 <= "0010"; -- 24
    when "00011001" => d1 <= "0101"; d2 <= "0010"; -- 25
    when "00011010" => d1 <= "0110"; d2 <= "0010"; -- 26
    when "00011011" => d1 <= "0111"; d2 <= "0010"; -- 27
    when "00011100" => d1 <= "1000"; d2 <= "0010"; -- 28
    when "00011101" => d1 <= "1001"; d2 <= "0010"; -- 29
    when "00011110" => d1 <= "0000"; d2 <= "0011"; -- 30
    when "00011111" => d1 <= "0001"; d2 <= "0011"; -- 31
    when "00100000" => d1 <= "0010"; d2 <= "0011"; -- 32
    when "00100001" => d1 <= "0011"; d2 <= "0011"; -- 33
    when "00100010" => d1 <= "0100"; d2 <= "0011"; -- 34
    when "00100011" => d1 <= "0101"; d2 <= "0011"; -- 35
    when "00100100" => d1 <= "0110"; d2 <= "0011"; -- 36
    when "00100101" => d1 <= "0111"; d2 <= "0011"; -- 37
    when "00100110" => d1 <= "1000"; d2 <= "0011"; -- 38
    when "00100111" => d1 <= "1001"; d2 <= "0011"; -- 39
    when "00101000" => d1 <= "0000"; d2 <= "0100"; -- 40
    when "00101001" => d1 <= "0001"; d2 <= "0100"; -- 41
    when "00101010" => d1 <= "0010"; d2 <= "0100"; -- 42
    when "00101011" => d1 <= "0011"; d2 <= "0100"; -- 43
    when "00101100" => d1 <= "0100"; d2 <= "0100"; -- 44
    when "00101101" => d1 <= "0101"; d2 <= "0100"; -- 45
    when "00101110" => d1 <= "0110"; d2 <= "0100"; -- 46
    when "00101111" => d1 <= "0111"; d2 <= "0100"; -- 47
    when "00110000" => d1 <= "1000"; d2 <= "0100"; -- 48
    when "00110001" => d1 <= "1001"; d2 <= "0100"; -- 49
    when "00110010" => d1 <= "0000"; d2 <= "0101"; -- 50
    when "00110011" => d1 <= "0001"; d2 <= "0101"; -- 51
    when "00110100" => d1 <= "0010"; d2 <= "0101"; -- 52
    when "00110101" => d1 <= "0011"; d2 <= "0101"; -- 53
    when "00110110" => d1 <= "0100"; d2 <= "0101"; -- 54
    when "00110111" => d1 <= "0101"; d2 <= "0101"; -- 55
    when "00111000" => d1 <= "0110"; d2 <= "0101"; -- 56
    when "00111001" => d1 <= "0111"; d2 <= "0101"; -- 57
    when "00111010" => d1 <= "1000"; d2 <= "0101"; -- 58
    when "00111011" => d1 <= "1001"; d2 <= "0101"; -- 59
	 when "00111100" => d1 <= "0000"; d2 <= "0110"; -- 60
    when "00111101" => d1 <= "0001"; d2 <= "0110"; -- 61
    when "00111110" => d1 <= "0010"; d2 <= "0110"; -- 62
    when "00111111" => d1 <= "0011"; d2 <= "0110"; -- 63
    when "01000000" => d1 <= "0100"; d2 <= "0110"; -- 64
    when "01000001" => d1 <= "0101"; d2 <= "0110"; -- 65
    when "01000010" => d1 <= "0110"; d2 <= "0110"; -- 66
    when "01000011" => d1 <= "0111"; d2 <= "0110"; -- 67
    when "01000100" => d1 <= "1000"; d2 <= "0110"; -- 68
    when "01000101" => d1 <= "1001"; d2 <= "0110"; -- 69
    when "01000110" => d1 <= "0000"; d2 <= "0111"; -- 70
    when "01000111" => d1 <= "0001"; d2 <= "0111"; -- 71
    when "01001000" => d1 <= "0010"; d2 <= "0111"; -- 72
    when "01001001" => d1 <= "0011"; d2 <= "0111"; -- 73
    when "01001010" => d1 <= "0100"; d2 <= "0111"; -- 74
    when "01001011" => d1 <= "0101"; d2 <= "0111"; -- 75
    when "01001100" => d1 <= "0110"; d2 <= "0111"; -- 76
    when "01001101" => d1 <= "0111"; d2 <= "0111"; -- 77
    when "01001110" => d1 <= "1000"; d2 <= "0111"; -- 78
    when "01001111" => d1 <= "1001"; d2 <= "0111"; -- 79
    when "01010000" => d1 <= "0000"; d2 <= "1000"; -- 80
    when "01010001" => d1 <= "0001"; d2 <= "1000"; -- 81
    when "01010010" => d1 <= "0010"; d2 <= "1000"; -- 82
    when "01010011" => d1 <= "0011"; d2 <= "1000"; -- 83
    when "01010100" => d1 <= "0100"; d2 <= "1000"; -- 84
    when "01010101" => d1 <= "0101"; d2 <= "1000"; -- 85
    when "01010110" => d1 <= "0110"; d2 <= "1000"; -- 86
    when "01010111" => d1 <= "0111"; d2 <= "1000"; -- 87
    when "01011000" => d1 <= "1000"; d2 <= "1000"; -- 88
    when "01011001" => d1 <= "1001"; d2 <= "1000"; -- 89
    when "01011010" => d1 <= "0000"; d2 <= "1001"; -- 90
    when "01011011" => d1 <= "0001"; d2 <= "1001"; -- 91
    when "01011100" => d1 <= "0010"; d2 <= "1001"; -- 92
    when "01011101" => d1 <= "0011"; d2 <= "1001"; -- 93
    when "01011110" => d1 <= "0100"; d2 <= "1001"; -- 94
    when "01011111" => d1 <= "0101"; d2 <= "1001"; -- 95
    when "01100000" => d1 <= "0110"; d2 <= "1001"; -- 96
    when "01100001" => d1 <= "0111"; d2 <= "1001"; -- 97
    when "01100010" => d1 <= "1000"; d2 <= "1001"; -- 98
    when "01100011" => d1 <= "1001"; d2 <= "1001"; -- 99
    when others =>
        d1 <= "0000"; d2 <= "0000";
end case;
					
					
				
		end process;

end architecture;